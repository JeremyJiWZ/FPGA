`timescale 1ns / 1ps
module Anti_jitter(input wire clk, 
						 input wire [3:0] button,
						 input wire [7:0] SW, 
						 output reg [3:0]button_out,
						 output reg [3:0]button_pulse,
						 output reg [7:0] SW_OK,
						 output reg rst

						);
	 
endmodule
